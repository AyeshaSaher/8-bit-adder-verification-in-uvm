interface adder_if(input logic clk);
  logic [7:0] operand_a;
  logic [7:0] operand_b;
  logic [7:0] sum;
endinterface
